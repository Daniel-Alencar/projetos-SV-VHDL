module hello;

    initial $display("Hello, FPGA!");
    
endmodule
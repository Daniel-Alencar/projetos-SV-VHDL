module porta_and (
  input A, B,
  output X
);
  assign X = A & B;
endmodule